`timescale 1ns / 1ps

module cbrt (
	input clk_i,
	input rst_i ,
	input [7 : 0] a_bi,
	output busy_o,
	output reg [3 : 0] y_bo
);

	localparam IDLE = 3'b000;
	localparam STATE1 = 3'b001;
	localparam STATE2 = 3'b010;
	localparam STATE3 = 3'b011;
	localparam STATE4 = 3'b100;
	localparam STATE5 = 3'b101;
	localparam STATE6 = 3'b110;
	localparam STATE7 = 3'b111;

	reg [7 : 0] a;

	reg [3 : 0] r, m;
	reg [7 : 0] n, p;

	reg [2 : 0] state;
	reg [2 : 0] state_next;

	reg [7:0] mult2_i1;
    reg [7:0] mult2_i2;
    wire [15:0] mult2_out;
    reg mult2_reset;
    wire mult2_busy;

    mult mult2(
        .clk_i(clk_i),
        .rst_i(mult2_reset),
        .a_bi(mult2_i1),
        .b_bi(mult2_i2),
        .busy_o(mult2_busy),
        .y_bo(mult2_out)
    );

	assign busy_o = rst_i | (state != 0);
	
	always @(posedge clk_i) 
        if (rst_i) begin
            state <= STATE1;
        end else begin
            state <= state_next;
        end

    always @* begin
        case(state)
            IDLE: state_next = IDLE;
            STATE1: state_next = (m != 0) ? STATE2 : IDLE;
            STATE2: state_next = mult2_busy ? STATE2 : STATE3;
            STATE3: state_next = mult2_busy ? STATE3 : STATE4;
            STATE4: state_next = STATE1;
        endcase
    end

    always @(posedge clk_i) begin
        if (rst_i) begin
            a <= a_bi;
            p <= 0;
            r <= 4;
            m <= 4;
            y_bo <= 0;
            mult2_reset <= 0;
        end else begin
	        case (state)
	            IDLE:
	                begin
                        y_bo <= r << 1;
                        if(p==1) begin
                            y_bo <= (r-1)<<1;
                        end
	                end
	            STATE1:
	                begin
	                   y_bo <= r;
	                   if (|m) begin
	                       mult2_reset <= 1;
	                       mult2_i1 <= r;
	                       mult2_i2 <= r;
	                   end
	                end
	            STATE2:
	                begin
	                    if (mult2_busy) begin
	                        mult2_reset <= 0;
	                    end else begin
	                        mult2_reset <= 1;
	                        mult2_i1 <= mult2_out;
	                        mult2_i2 <= r;
	                    end
	                end
	            STATE3:
	                begin
	                    mult2_reset <= 0;
	                    if (!mult2_busy) begin
	                        if (a == mult2_out) begin
	                            m <= 0;
	                        end else if (a < mult2_out) begin
	                            r <= r - m;
	                        end else begin
	                            r <= r + m;
	                        end
                            if(a<125) 
                                begin 
                                    if(a>64) begin
                                        p<=1; end
                                end
                                
                            if(a<27) 
                                begin 
                                    if(a>8) begin
                                        p<=1; end
                                end
	                    end
	                end
	            STATE4:
	                begin
	                    if (m >= 1) begin
	                        m <= m >> 1;
	                    end
	                 end
	        endcase
        end
    end
endmodule